library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY MEMORY IS
	PORT( ADDRESS: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		ENABLE, SAMPLE: IN STD_LOGIC; -- sample is the timed signal form FSM
		DATAOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
		
	END MEMORY;
	ARCHITECTURE RAM OF MEMORY IS
		TYPE WAVE IS ARRAY (0 TO 1023) OF STD_LOGIC_VECTOR(7 DOWNTO 0); -- Array storing sample values.
		--First two bits in address represent wave type. 00 is sine, 01 square, 10 triangle, and 11 sawtooth. Max sample number is 256 for each type.
		--This was originally implemented as a 2D array but was changed during debugging. It could still be implemented as such to make it easier to
		--replace types with different ones but we'll leave it as such due to project time restraints.
		CONSTANT SAMPLEVALUE : WAVE := ("10000000", "10000011", "10000110", "10001001", "10001100", "10001111", "10010010", "10010101", "10011000",
		"10011011", "10011110", "10100010", "10100101", "10100111", "10101010", "10101101", "10110000", "10110011", "10110110", "10111001", "10111100",
		"10111110", "11000001", "11000100", "11000110", "11001001", "11001011", "11001110", "11010000", "11010011", "11010101", "11010111", "11011010",
		"11011100", "11011110", "11100000", "11100010", "11100100", "11100110", "11101000", "11101010", "11101011", "11101101", "11101110", "11110000",
		"11110001", "11110011", "11110100", "11110101", "11110110", "11111000", "11111001", "11111010", "11111010", "11111011", "11111100", "11111101",
		"11111101", "11111110", "11111110", "11111110", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111110",
		"11111110", "11111110", "11111101", "11111101", "11111100", "11111011", "11111010", "11111010", "11111001", "11111000", "11110110", "11110101",
		"11110100", "11110011", "11110001", "11110000", "11101110", "11101101", "11101011", "11101010", "11101000", "11100110", "11100100", "11100010",
		"11100000", "11011110", "11011100", "11011010", "11010111", "11010101", "11010011", "11010000", "11001110", "11001011", "11001001", "11000110",
		"11000100", "11000001", "10111110", "10111100", "10111001", "10110110", "10110011", "10110000", "10101101", "10101010", "10100111", "10100101",
		"10100010", "10011110", "10011011", "10011000", "10010101", "10010010", "10001111", "10001100", "10001001", "10000110", "10000011", "10000000",
		"01111100", "01111001", "01110110", "01110011", "01110000", "01101101", "01101010", "01100111", "01100100", "01100001", "01011101", "01011010",
		"01011000", "01010101", "01010010", "01001111", "01001100", "01001001", "01000110", "01000011", "01000001", "00111110", "00111011", "00111001",
		"00110110", "00110100", "00110001", "00101111", "00101100", "00101010", "00101000", "00100101", "00100011", "00100001", "00011111", "00011101",
		"00011011", "00011001", "00010111", "00010101", "00010100", "00010010", "00010001", "00001111", "00001110", "00001100", "00001011", "00001010",
		"00001001", "00000111", "00000110", "00000101", "00000101", "00000100", "00000011", "00000010", "00000010", "00000001", "00000001", "00000001",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000001", "00000001", "00000001", "00000010", "00000010",
		"00000011", "00000100", "00000101", "00000101", "00000110", "00000111", "00001001", "00001010", "00001011", "00001100", "00001110", "00001111",
		"00010001", "00010010", "00010100", "00010101", "00010111", "00011001", "00011011", "00011101", "00011111", "00100001", "00100011", "00100101",
		"00101000", "00101010", "00101100", "00101111", "00110001", "00110100", "00110110", "00111001", "00111011", "00111110", "01000001", "01000011",
		"01000110", "01001001", "01001100", "01001111", "01010010", "01010101", "01011000", "01011010", "01011101", "01100001", "01100100", "01100111",
		"01101010", "01101101", "01110000", "01110011", "01110110", "01111001", "01111100",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
		"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111",
		"11111111", "11111111", "11111111", "11111111",
		"00000000", "00000010", "00000100", "00000110", "00001000", "00001010", "00001100", "00001110", "00010000", "00010010", "00010100", "00010110",
 		"00011000", "00011010", "00011100", "00011110", "00100000", "00100010", "00100100", "00100110", "00101000", "00101010", "00101100", "00101110",
		"00110000", "00110010", "00110100", "00110110", "00111000", "00111010", "00111100", "00111110", "01000000", "01000010", "01000100", "01000110",
		"01001000", "01001010", "01001100", "01001110", "01010000", "01010010", "01010100", "01010110", "01011000", "01011010", "01011100", "01011110", 
		"01100000", "01100010", "01100100", "01100110", "01101000", "01101010", "01101100", "01101110", "01110000", "01110010", "01110100", "01110110", 
		"01111000", "01111010", "01111100", "01111110", "10000000", "10000001", "10000011", "10000101", "10000111", "10001001", "10001011", "10001101", 
		"10001111", "10010001", "10010011", "10010101", "10010111", "10011001", "10011011", "10011101", "10011111", "10100001", "10100011", "10100101", 
		"10100111", "10101001", "10101011", "10101101", "10101111", "10110001", "10110011", "10110101", "10110111", "10111001", "10111011", "10111101", 
		"10111111", "11000001", "11000011", "11000101", "11000111", "11001001", "11001011", "11001101", "11001111", "11010001", "11010011", "11010101", 
		"11010111", "11011001", "11011011", "11011101", "11011111", "11100001", "11100011", "11100101", "11100111", "11101001", "11101011", "11101101", 
		"11101111", "11110001", "11110011", "11110101", "11110111", "11111001", "11111011", "11111101", "11111111", "11111101", "11111011", "11111001", 
		"11110111", "11110101", "11110011", "11110001", "11101111", "11101101", "11101011", "11101001", "11100111", "11100101", "11100011", "11100001", 
		"11011111", "11011101", "11011011", "11011001", "11010111", "11010101", "11010011", "11010001", "11001111", "11001101", "11001011", "11001001", 
		"11000111", "11000101", "11000011", "11000001", "10111111", "10111101", "10111011", "10111001", "10110111", "10110101", "10110011", "10110001", 
		"10101111", "10101101", "10101011", "10101001", "10100111", "10100101", "10100011", "10100001", "10011111", "10011101", "10011011", "10011001", 
		"10010111", "10010101", "10010011", "10010001", "10001111", "10001101", "10001011", "10001001", "10000111", "10000101", "10000011", "10000001", 
		"10000000", "01111110", "01111100", "01111010", "01111000", "01110110", "01110100", "01110010", "01110000", "01101110", "01101100", "01101010", 
		"01101000", "01100110", "01100100", "01100010", "01100000", "01011110", "01011100", "01011010", "01011000", "01010110", "01010100", "01010010", 
		"01010000", "01001110", "01001100", "01001010", "01001000", "01000110", "01000100", "01000010", "01000000", "00111110", "00111100", "00111010", 
		"00111000", "00110110", "00110100", "00110010", "00110000", "00101110", "00101100", "00101010", "00101000", "00100110", "00100100", "00100010", 
		"00100000", "00011110", "00011100", "00011010", "00011000", "00010110", "00010100", "00010010", "00010000", "00001110", "00001100", "00001010", 
		"00001000", "00000110", "00000100", "00000010",
		"00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111", "00001000", "00001001", "00001010", "00001011",
		"00001100", "00001101", "00001110", "00001111", "00010000", "00010001", "00010010", "00010011", "00010100", "00010101", "00010110", "00010111",
		"00011000", "00011001", "00011010", "00011011", "00011100", "00011101", "00011110", "00011111", "00100000", "00100001", "00100010", "00100011",
		"00100100", "00100101", "00100110", "00100111", "00101000", "00101001", "00101010", "00101011", "00101100", "00101101", "00101110", "00101111",
		"00110000", "00110001", "00110010", "00110011", "00110100", "00110101", "00110110", "00110111", "00111000", "00111001", "00111010", "00111011",
		"00111100", "00111101", "00111110", "00111111", "01000000", "01000001", "01000010", "01000011", "01000100", "01000101", "01000110", "01000111",
		"01001000", "01001001", "01001010", "01001011", "01001100", "01001101", "01001110", "01001111", "01010000", "01010001", "01010010", "01010011",
		"01010100", "01010101", "01010110", "01010111", "01011000", "01011001", "01011010", "01011011", "01011100", "01011101", "01011110", "01011111",
		"01100000", "01100001", "01100010", "01100011", "01100100", "01100101", "01100110", "01100111", "01101000", "01101001", "01101010", "01101011",
		"01101100", "01101101", "01101110", "01101111", "01110000", "01110001", "01110010", "01110011", "01110100", "01110101", "01110110", "01110111",
		"01111000", "01111001", "01111010", "01111011", "01111100", "01111101", "01111110", "01111111", "10000000", "10000001", "10000010", "10000011",
		"10000100", "10000101", "10000110", "10000111", "10001000", "10001001", "10001010", "10001011", "10001100", "10001101", "10001110", "10001111",
		"10010000", "10010001", "10010010", "10010011", "10010100", "10010101", "10010110", "10010111", "10011000", "10011001", "10011010", "10011011",
		"10011100", "10011101", "10011110", "10011111", "10100000", "10100001", "10100010", "10100011", "10100100", "10100101", "10100110", "10100111",
		"10101000", "10101001", "10101010", "10101011", "10101100", "10101101", "10101110", "10101111", "10110000", "10110001", "10110010", "10110011",
		"10110100", "10110101", "10110110", "10110111", "10111000", "10111001", "10111010", "10111011", "10111100", "10111101", "10111110", "10111111",
		"11000000", "11000001", "11000010", "11000011", "11000100", "11000101", "11000110", "11000111", "11001000", "11001001", "11001010", "11001011",
		"11001100", "11001101", "11001110", "11001111", "11010000", "11010001", "11010010", "11010011", "11010100", "11010101", "11010110", "11010111",
		"11011000", "11011001", "11011010", "11011011", "11011100", "11011101", "11011110", "11011111", "11100000", "11100001", "11100010", "11100011",
		"11100100", "11100101", "11100110", "11100111", "11101000", "11101001", "11101010", "11101011", "11101100", "11101101", "11101110", "11101111",
		"11110000", "11110001", "11110010", "11110011", "11110100", "11110101", "11110110", "11110111", "11111000", "11111001", "11111010", "11111011",
		"11111100", "11111101", "11111110", "11111111"
		);
		
		
		SIGNAL TTEMP : STD_LOGIC_VECTOR(7 DOWNTO 0);
		BEGIN
		PROCESS(ADDRESS, ENABLE, SAMPLE)
		BEGIN
			IF((ENABLE and SAMPLE) = '1')THEN
				TTEMP <= SAMPLEVALUE(TO_INTEGER(UNSIGNED(ADDRESS(9 DOWNTO 0))));
				ELSE
				TTEMP <= TTEMP;
			END IF;
		END PROCESS;
		DATAOUT <= TTEMP;
	END RAM;