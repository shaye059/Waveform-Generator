library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY WAVEFORM_TOP IS
	PORT(
		WAVE_TYPE: IN STD_LOGIC_VECTOR(1 DOWNTO 0); 	-- CH_WF
		PERIOD: IN STD_LOGIC_VECTOR(9 DOWNTO 0); 	--CH_P
		SAMPLE_RATE: IN STD_LOGIC_VECTOR(7 DOWNTO 0); 	--CH_SR
		START: IN STD_LOGIC; 				--START SIGNAL
		CLOCK : IN STD_LOGIC; 				--SYSTEM CLOCK
		RESET : IN STD_LOGIC;				--RESTART
		DATA_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);

END WAVEFORM_TOP;

ARCHITECTURE TOP_STRU OF WAVEFORM_TOP IS
	SIGNAL P: STD_LOGIC_VECTOR(9 DOWNTO 0);
	SIGNAL CC: STD_LOGIC;
	SIGNAL R: STD_LOGIC;
	SIGNAL FULL: STD_LOGIC;
	SIGNAL CS: STD_LOGIC;
	SIGNAL EN: STD_LOGIC;
	SIGNAL LP: STD_LOGIC;
	SIGNAL ADDR: STD_LOGIC_VECTOR(9 DOWNTO 0);
	SIGNAL DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);

	COMPONENT FSM_CTRL
		PORT (CLK	:	IN STD_LOGIC;
		RST	:	IN STD_LOGIC;
		ST	:	IN STD_LOGIC;
		CH_WF	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		CH_P	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		CH_SR	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		FULL	:	IN STD_LOGIC;

		P		:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		CC		:	OUT STD_LOGIC;
		CS		:	OUT STD_LOGIC;
		EN		:	OUT STD_LOGIC;
		LP		:	OUT STD_LOGIC;
		R		:	OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT COUNTER
		PORT(CC : IN STD_LOGIC;
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		P : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		ADDR : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
		FULL : OUT STD_LOGIC
		);
	END COMPONENT;

	COMPONENT MEMORY
		PORT( ADDRESS: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		ENABLE, SAMPLE: IN STD_LOGIC; -- sample is the timed signal form FSM
		DATAOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT DATA_LATCH_LOGIC
		PORT(D_IN		: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		LP		: IN STD_LOGIC;
		D_OUT		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		);
	END COMPONENT;

BEGIN
	L1: FSM_CTRL PORT MAP (CLOCK, RESET, START, WAVE_TYPE, PERIOD, SAMPLE_RATE, FULL, P, CC, CS, EN, LP, R);
	L2: COUNTER PORT MAP (CC, CLOCK, R, P, ADDR, FULL);
	L3: MEMORY PORT MAP (ADDR, EN, CS, DATA);
	L4: DATA_LATCH_LOGIC PORT MAP (DATA, LP, DATA_OUT);

END TOP_STRU;

